library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;



package waveform_lut is

signal i : integer range 0 to 127:= 0;
signal j : integer range 0 to 127:=0;
signal k : integer range 0 to 127:=0;

type sin_lut is array (0 to 127) of integer; 
 
constant S_LUT : sin_lut  := ( 
0 => 512 , 
1 => 537 , 
2 => 562 , 
3 => 587 , 
4 => 611 , 
5 => 636 , 
6 => 660 , 
7 => 684 , 
8 => 707 , 
9 => 730 , 
10 => 753 , 
11 => 774 , 
12 => 796 , 
13 => 816 , 
14 => 836 , 
15 => 855 , 
16 => 873 , 
17 => 890 , 
18 => 907 , 
19 => 922 , 
20 => 937 , 
21 => 950 , 
22 => 962 , 
23 => 974 , 
24 => 984 , 
25 => 993 , 
26 => 1001 , 
27 => 1008 , 
28 => 1013 , 
29 => 1017 , 
30 => 1020 , 
31 => 1022 , 
32 => 1022 , 
33 => 1020 , 
34 => 1017 , 
35 => 1013 , 
36 => 1008 , 
37 => 1001 , 
38 => 993 , 
39 => 984 , 
40 => 974 , 
41 => 962 , 
42 => 950 , 
43 => 937 , 
44 => 922 , 
45 => 907 , 
46 => 890 , 
47 => 873 , 
48 => 855 , 
49 => 836 , 
50 => 816 , 
51 => 796 , 
52 => 774 , 
53 => 753 , 
54 => 730 , 
55 => 707 , 
56 => 684 , 
57 => 660 , 
58 => 636 , 
59 => 611 , 
60 => 587 , 
61 => 562 , 
62 => 537 , 
63 => 512 , 
64 => 512 , 
65 => 487 , 
66 => 462 , 
67 => 437 , 
68 => 413 , 
69 => 388 , 
70 => 364 , 
71 => 340 , 
72 => 317 , 
73 => 294 , 
74 => 271 , 
75 => 250 , 
76 => 228 , 
77 => 208 , 
78 => 188 , 
79 => 169 , 
80 => 151 , 
81 => 134 , 
82 => 117 , 
83 => 102 , 
84 => 87 , 
85 => 74 , 
86 => 62 , 
87 => 50 , 
88 => 40 , 
89 => 31 , 
90 => 23 , 
91 => 16 , 
92 => 11 , 
93 => 7 , 
94 => 4 , 
95 => 2 , 
96 => 2 , 
97 => 4 , 
98 => 7 , 
99 => 11 , 
100 => 16 , 
101 => 23 , 
102 => 31 , 
103 => 40 , 
104 => 50 , 
105 => 62 , 
106 => 74 , 
107 => 87 , 
108 => 102 , 
109 => 117 , 
110 => 134 , 
111 => 151 , 
112 => 169 , 
113 => 188 , 
114 => 208 , 
115 => 228 , 
116 => 250 , 
117 => 271 , 
118 => 294 , 
119 => 317 , 
120 => 340 , 
121 => 364 , 
122 => 388 , 
123 => 413 , 
124 => 437 , 
125 => 462 , 
126 => 487 , 
127 => 512  
);

type tri_lut is array (0 to 511) of integer; 
 
constant T_LUT : tri_lut  := ( 
0 => 512 , 
1 => 516 , 
2 => 520 , 
3 => 524 , 
4 => 528 , 
5 => 532 , 
6 => 536 , 
7 => 540 , 
8 => 544 , 
9 => 548 , 
10 => 552 , 
11 => 556 , 
12 => 560 , 
13 => 564 , 
14 => 568 , 
15 => 572 , 
16 => 576 , 
17 => 580 , 
18 => 584 , 
19 => 588 , 
20 => 592 , 
21 => 596 , 
22 => 600 , 
23 => 604 , 
24 => 608 , 
25 => 612 , 
26 => 616 , 
27 => 620 , 
28 => 624 , 
29 => 628 , 
30 => 632 , 
31 => 636 , 
32 => 640 , 
33 => 644 , 
34 => 648 , 
35 => 652 , 
36 => 656 , 
37 => 661 , 
38 => 665 , 
39 => 669 , 
40 => 673 , 
41 => 677 , 
42 => 681 , 
43 => 685 , 
44 => 689 , 
45 => 693 , 
46 => 697 , 
47 => 701 , 
48 => 705 , 
49 => 709 , 
50 => 713 , 
51 => 717 , 
52 => 721 , 
53 => 725 , 
54 => 729 , 
55 => 733 , 
56 => 737 , 
57 => 741 , 
58 => 745 , 
59 => 749 , 
60 => 753 , 
61 => 757 , 
62 => 761 , 
63 => 765 , 
64 => 769 , 
65 => 773 , 
66 => 777 , 
67 => 781 , 
68 => 785 , 
69 => 789 , 
70 => 793 , 
71 => 797 , 
72 => 801 , 
73 => 806 , 
74 => 810 , 
75 => 814 , 
76 => 818 , 
77 => 822 , 
78 => 826 , 
79 => 830 , 
80 => 834 , 
81 => 838 , 
82 => 842 , 
83 => 846 , 
84 => 850 , 
85 => 854 , 
86 => 858 , 
87 => 862 , 
88 => 866 , 
89 => 870 , 
90 => 874 , 
91 => 878 , 
92 => 882 , 
93 => 886 , 
94 => 890 , 
95 => 894 , 
96 => 898 , 
97 => 902 , 
98 => 906 , 
99 => 910 , 
100 => 914 , 
101 => 918 , 
102 => 922 , 
103 => 926 , 
104 => 930 , 
105 => 934 , 
106 => 938 , 
107 => 942 , 
108 => 946 , 
109 => 951 , 
110 => 955 , 
111 => 959 , 
112 => 963 , 
113 => 967 , 
114 => 971 , 
115 => 975 , 
116 => 979 , 
117 => 983 , 
118 => 987 , 
119 => 991 , 
120 => 995 , 
121 => 999 , 
122 => 1003 , 
123 => 1007 , 
124 => 1011 , 
125 => 1015 , 
126 => 1019 , 
127 => 1023 , 
128 => 1023 , 
129 => 1019 , 
130 => 1015 , 
131 => 1011 , 
132 => 1007 , 
133 => 1003 , 
134 => 999 , 
135 => 995 , 
136 => 991 , 
137 => 987 , 
138 => 983 , 
139 => 979 , 
140 => 975 , 
141 => 971 , 
142 => 967 , 
143 => 963 , 
144 => 959 , 
145 => 955 , 
146 => 951 , 
147 => 946 , 
148 => 942 , 
149 => 938 , 
150 => 934 , 
151 => 930 , 
152 => 926 , 
153 => 922 , 
154 => 918 , 
155 => 914 , 
156 => 910 , 
157 => 906 , 
158 => 902 , 
159 => 898 , 
160 => 894 , 
161 => 890 , 
162 => 886 , 
163 => 882 , 
164 => 878 , 
165 => 874 , 
166 => 870 , 
167 => 866 , 
168 => 862 , 
169 => 858 , 
170 => 854 , 
171 => 850 , 
172 => 846 , 
173 => 842 , 
174 => 838 , 
175 => 834 , 
176 => 830 , 
177 => 826 , 
178 => 822 , 
179 => 818 , 
180 => 814 , 
181 => 810 , 
182 => 806 , 
183 => 801 , 
184 => 797 , 
185 => 793 , 
186 => 789 , 
187 => 785 , 
188 => 781 , 
189 => 777 , 
190 => 773 , 
191 => 769 , 
192 => 765 , 
193 => 761 , 
194 => 757 , 
195 => 753 , 
196 => 749 , 
197 => 745 , 
198 => 741 , 
199 => 737 , 
200 => 733 , 
201 => 729 , 
202 => 725 , 
203 => 721 , 
204 => 717 , 
205 => 713 , 
206 => 709 , 
207 => 705 , 
208 => 701 , 
209 => 697 , 
210 => 693 , 
211 => 689 , 
212 => 685 , 
213 => 681 , 
214 => 677 , 
215 => 673 , 
216 => 669 , 
217 => 665 , 
218 => 661 , 
219 => 656 , 
220 => 652 , 
221 => 648 , 
222 => 644 , 
223 => 640 , 
224 => 636 , 
225 => 632 , 
226 => 628 , 
227 => 624 , 
228 => 620 , 
229 => 616 , 
230 => 612 , 
231 => 608 , 
232 => 604 , 
233 => 600 , 
234 => 596 , 
235 => 592 , 
236 => 588 , 
237 => 584 , 
238 => 580 , 
239 => 576 , 
240 => 572 , 
241 => 568 , 
242 => 564 , 
243 => 560 , 
244 => 556 , 
245 => 552 , 
246 => 548 , 
247 => 544 , 
248 => 540 , 
249 => 536 , 
250 => 532 , 
251 => 528 , 
252 => 524 , 
253 => 520 , 
254 => 516 , 
255 => 512 , 
256 => 511 , 
257 => 507 , 
258 => 503 , 
259 => 499 , 
260 => 495 , 
261 => 491 , 
262 => 487 , 
263 => 483 , 
264 => 479 , 
265 => 475 , 
266 => 471 , 
267 => 467 , 
268 => 463 , 
269 => 459 , 
270 => 455 , 
271 => 451 , 
272 => 447 , 
273 => 443 , 
274 => 439 , 
275 => 434 , 
276 => 430 , 
277 => 426 , 
278 => 422 , 
279 => 418 , 
280 => 414 , 
281 => 410 , 
282 => 406 , 
283 => 402 , 
284 => 398 , 
285 => 394 , 
286 => 390 , 
287 => 386 , 
288 => 382 , 
289 => 378 , 
290 => 374 , 
291 => 370 , 
292 => 366 , 
293 => 362 , 
294 => 358 , 
295 => 354 , 
296 => 350 , 
297 => 346 , 
298 => 342 , 
299 => 338 , 
300 => 334 , 
301 => 330 , 
302 => 326 , 
303 => 322 , 
304 => 318 , 
305 => 314 , 
306 => 310 , 
307 => 306 , 
308 => 302 , 
309 => 298 , 
310 => 294 , 
311 => 289 , 
312 => 285 , 
313 => 281 , 
314 => 277 , 
315 => 273 , 
316 => 269 , 
317 => 265 , 
318 => 261 , 
319 => 257 , 
320 => 253 , 
321 => 249 , 
322 => 245 , 
323 => 241 , 
324 => 237 , 
325 => 233 , 
326 => 229 , 
327 => 225 , 
328 => 221 , 
329 => 217 , 
330 => 213 , 
331 => 209 , 
332 => 205 , 
333 => 201 , 
334 => 197 , 
335 => 193 , 
336 => 189 , 
337 => 185 , 
338 => 181 , 
339 => 177 , 
340 => 173 , 
341 => 169 , 
342 => 165 , 
343 => 161 , 
344 => 157 , 
345 => 153 , 
346 => 149 , 
347 => 144 , 
348 => 140 , 
349 => 136 , 
350 => 132 , 
351 => 128 , 
352 => 124 , 
353 => 120 , 
354 => 116 , 
355 => 112 , 
356 => 108 , 
357 => 104 , 
358 => 100 , 
359 => 96 , 
360 => 92 , 
361 => 88 , 
362 => 84 , 
363 => 80 , 
364 => 76 , 
365 => 72 , 
366 => 68 , 
367 => 64 , 
368 => 60 , 
369 => 56 , 
370 => 52 , 
371 => 48 , 
372 => 44 , 
373 => 40 , 
374 => 36 , 
375 => 32 , 
376 => 28 , 
377 => 24 , 
378 => 20 , 
379 => 16 , 
380 => 12 , 
381 => 8 , 
382 => 4 , 
383 => 0 , 
384 => 0 , 
385 => 4 , 
386 => 8 , 
387 => 12 , 
388 => 16 , 
389 => 20 , 
390 => 24 , 
391 => 28 , 
392 => 32 , 
393 => 36 , 
394 => 40 , 
395 => 44 , 
396 => 48 , 
397 => 52 , 
398 => 56 , 
399 => 60 , 
400 => 64 , 
401 => 68 , 
402 => 72 , 
403 => 76 , 
404 => 80 , 
405 => 84 , 
406 => 88 , 
407 => 92 , 
408 => 96 , 
409 => 100 , 
410 => 104 , 
411 => 108 , 
412 => 112 , 
413 => 116 , 
414 => 120 , 
415 => 124 , 
416 => 128 , 
417 => 132 , 
418 => 136 , 
419 => 140 , 
420 => 144 , 
421 => 149 , 
422 => 153 , 
423 => 157 , 
424 => 161 , 
425 => 165 , 
426 => 169 , 
427 => 173 , 
428 => 177 , 
429 => 181 , 
430 => 185 , 
431 => 189 , 
432 => 193 , 
433 => 197 , 
434 => 201 , 
435 => 205 , 
436 => 209 , 
437 => 213 , 
438 => 217 , 
439 => 221 , 
440 => 225 , 
441 => 229 , 
442 => 233 , 
443 => 237 , 
444 => 241 , 
445 => 245 , 
446 => 249 , 
447 => 253 , 
448 => 257 , 
449 => 261 , 
450 => 265 , 
451 => 269 , 
452 => 273 , 
453 => 277 , 
454 => 281 , 
455 => 285 , 
456 => 289 , 
457 => 294 , 
458 => 298 , 
459 => 302 , 
460 => 306 , 
461 => 310 , 
462 => 314 , 
463 => 318 , 
464 => 322 , 
465 => 326 , 
466 => 330 , 
467 => 334 , 
468 => 338 , 
469 => 342 , 
470 => 346 , 
471 => 350 , 
472 => 354 , 
473 => 358 , 
474 => 362 , 
475 => 366 , 
476 => 370 , 
477 => 374 , 
478 => 378 , 
479 => 382 , 
480 => 386 , 
481 => 390 , 
482 => 394 , 
483 => 398 , 
484 => 402 , 
485 => 406 , 
486 => 410 , 
487 => 414 , 
488 => 418 , 
489 => 422 , 
490 => 426 , 
491 => 430 , 
492 => 434 , 
493 => 439 , 
494 => 443 , 
495 => 447 , 
496 => 451 , 
497 => 455 , 
498 => 459 , 
499 => 463 , 
500 => 467 , 
501 => 471 , 
502 => 475 , 
503 => 479 , 
504 => 483 , 
505 => 487 , 
506 => 491 , 
507 => 495 , 
508 => 499 , 
509 => 503 , 
510 => 507 , 
511 => 511  
);




end waveform_lut;